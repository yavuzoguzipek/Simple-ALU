library verilog;
use verilog.vl_types.all;
entity MyXor is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end MyXor;
