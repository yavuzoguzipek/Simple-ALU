library verilog;
use verilog.vl_types.all;
entity demo is
end demo;
