library verilog;
use verilog.vl_types.all;
entity Sub4 is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end Sub4;
